`timescale 1ns / 1ps

module add_tb (
	
);
	
endmodule
